`timescale 1ns / 1ps

module testflow();

// Inputs

// Outputs

        
top UUT (/*
            .cnt_th(cnt_th),
            .dn_up(dn_up), 
            .timeout(timeout), 
            .cntout(cntout), 
            .n_reset(n_reset), 
            .enable(enable), 
            .clk(clk)*/
            );

 
endmodule