`timescale 1ns / 1ps
// Parameters:  SPI_MODE, can be 0, 1, 2, 3.
//              Can be configured in one of 4 modes:
//              Mode | Clock Polarity (CPOL/CKP) | Clock Phase (CPHA)
//               0   |             0             |        0
//               1   |             0             |        1
//               2   |             1             |        0
//               3   |             1             |        1
module spi_master(

    );
endmodule
