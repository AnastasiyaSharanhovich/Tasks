`timescale 1ns / 1ps

module apb_addr_dec(

    );
    
endmodule
