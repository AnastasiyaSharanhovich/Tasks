`timescale 1ns / 1ps
//sync_fifo
module fifo(

    );
endmodule
